library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity singen is
	PORT( 									
		angle: IN integer range 0 to 65535;
		sinAngle	:	OUT integer range 0 to 65535;
		cosAngle	:	OUT integer range 0 to 65535); -- 16 bit wide(0 to 2^[16-1])	
END singen;

ARCHITECTURE RTL OF singen IS
	type memory_type is array (0 to 4095) of integer range 0 to 65535;
	signal sine     :    memory_type :=(32768,32818,32868,32918,32969,33019,33069,33119,33170,33220,33270,33320,33371,33421,33471,33521,33572,33622,33672,33722,33773,33823,33873,33923,33974,34024,34074,34124,34175,34225,34275,34325,34375,34426,34476,34526,34576,34626,34677,34727,34777,34827,34877,34927,34978,35028,35078,35128,35178,35228,35278,35328,35379,35429,35479,35529,35579,35629,35679,35729,35779,35829,35879,35929,35979,36029,36079,36129,36179,36229,36279,36329,36379,36429,36479,36529,36579,36629,36679,36729,36779,36829,36878,36928,36978,37028,37078,37128,37177,37227,37277,37327,37377,37426,37476,37526,37576,37625,37675,37725,37774,37824,37874,37923,37973,38023,38072,38122,38171,38221,38271,38320,38370,38419,38469,38518,38568,38617,38666,38716,38765,38815,38864,38914,38963,39012,39062,39111,39160,39210,39259,39308,39357,39407,39456,39505,39554,39603,39652,39702,39751,39800,39849,39898,39947,39996,40045,40094,40143,40192,40241,40290,40339,40388,40437,40485,40534,40583,40632,40681,40729,40778,40827,40876,40924,40973,41022,41070,41119,41168,41216,41265,41313,41362,41410,41459,41507,41556,41604,41652,41701,41749,41797,41846,41894,41942,41991,42039,42087,42135,42183,42231,42280,42328,42376,42424,42472,42520,42568,42616,42664,42712,42759,42807,42855,42903,42951,42998,43046,43094,43142,43189,43237,43285,43332,43380,43427,43475,43522,43570,43617,43665,43712,43759,43807,43854,43901,43949,43996,44043,44090,44137,44184,44232,44279,44326,44373,44420,44467,44514,44561,44607,44654,44701,44748,44795,44841,44888,44935,44981,45028,45075,45121,45168,45214,45261,45307,45354,45400,45446,45493,45539,45585,45632,45678,45724,45770,45816,45862,45908,45954,46000,46046,46092,46138,46184,46230,46276,46322,46367,46413,46459,46504,46550,46596,46641,46687,46732,46778,46823,46868,46914,46959,47004,47050,47095,47140,47185,47230,47275,47320,47366,47410,47455,47500,47545,47590,47635,47680,47724,47769,47814,47858,47903,47948,47992,48037,48081,48125,48170,48214,48259,48303,48347,48391,48435,48480,48524,48568,48612,48656,48700,48744,48787,48831,48875,48919,48963,49006,49050,49093,49137,49181,49224,49267,49311,49354,49398,49441,49484,49527,49570,49614,49657,49700,49743,49786,49829,49872,49914,49957,50000,50043,50085,50128,50171,50213,50256,50298,50341,50383,50426,50468,50510,50552,50595,50637,50679,50721,50763,50805,50847,50889,50931,50972,51014,51056,51098,51139,51181,51222,51264,51305,51347,51388,51430,51471,51512,51553,51594,51636,51677,51718,51759,51800,51841,51881,51922,51963,52004,52044,52085,52126,52166,52207,52247,52287,52328,52368,52408,52449,52489,52529,52569,52609,52649,52689,52729,52769,52808,52848,52888,52927,52967,53007,53046,53086,53125,53164,53204,53243,53282,53321,53360,53399,53439,53477,53516,53555,53594,53633,53672,53710,53749,53788,53826,53865,53903,53941,53980,54018,54056,54094,54133,54171,54209,54247,54285,54323,54360,54398,54436,54474,54511,54549,54586,54624,54661,54699,54736,54773,54810,54848,54885,54922,54959,54996,55033,55069,55106,55143,55180,55216,55253,55289,55326,55362,55399,55435,55471,55508,55544,55580,55616,55652,55688,55724,55760,55795,55831,55867,55902,55938,55973,56009,56044,56080,56115,56150,56185,56221,56256,56291,56326,56361,56395,56430,56465,56500,56534,56569,56603,56638,56672,56707,56741,56775,56809,56843,56877,56912,56945,56979,57013,57047,57081,57114,57148,57182,57215,57248,57282,57315,57348,57382,57415,57448,57481,57514,57547,57580,57613,57645,57678,57711,57743,57776,57808,57841,57873,57905,57937,57969,58002,58034,58066,58098,58129,58161,58193,58225,58256,58288,58319,58351,58382,58413,58445,58476,58507,58538,58569,58600,58631,58662,58693,58723,58754,58784,58815,58845,58876,58906,58937,58967,58997,59027,59057,59087,59117,59147,59177,59206,59236,59266,59295,59325,59354,59383,59413,59442,59471,59500,59529,59558,59587,59616,59645,59673,59702,59731,59759,59788,59816,59844,59873,59901,59929,59957,59985,60013,60041,60069,60097,60124,60152,60179,60207,60234,60262,60289,60316,60344,60371,60398,60425,60452,60479,60505,60532,60559,60585,60612,60638,60665,60691,60717,60744,60770,60796,60822,60848,60874,60899,60925,60951,60976,61002,61027,61053,61078,61103,61129,61154,61179,61204,61229,61254,61279,61303,61328,61353,61377,61402,61426,61450,61475,61499,61523,61547,61571,61595,61619,61643,61666,61690,61714,61737,61761,61784,61807,61830,61854,61877,61900,61923,61946,61969,61991,62014,62037,62059,62082,62104,62127,62149,62171,62193,62215,62237,62259,62281,62303,62325,62346,62368,62389,62411,62432,62454,62475,62496,62517,62538,62559,62580,62601,62622,62642,62663,62683,62704,62724,62745,62765,62785,62805,62825,62845,62865,62885,62905,62924,62944,62964,62983,63003,63022,63041,63060,63080,63099,63118,63136,63155,63174,63193,63211,63230,63248,63267,63285,63303,63322,63340,63358,63376,63394,63412,63429,63447,63465,63482,63500,63517,63534,63552,63569,63586,63603,63620,63637,63654,63670,63687,63704,63720,63737,63753,63769,63786,63802,63818,63834,63850,63866,63882,63897,63913,63929,63944,63960,63975,63990,64005,64021,64036,64051,64066,64080,64095,64110,64125,64139,64154,64168,64182,64197,64211,64225,64239,64253,64267,64281,64294,64308,64322,64335,64349,64362,64375,64388,64402,64415,64428,64441,64453,64466,64479,64491,64504,64517,64529,64541,64553,64566,64578,64590,64602,64614,64625,64637,64649,64660,64672,64683,64695,64706,64717,64728,64739,64750,64761,64772,64783,64793,64804,64815,64825,64835,64846,64856,64866,64876,64886,64896,64906,64916,64925,64935,64944,64954,64963,64973,64982,64991,65000,65009,65018,65027,65036,65044,65053,65062,65070,65079,65087,65095,65103,65111,65119,65127,65135,65143,65151,65158,65166,65173,65181,65188,65195,65203,65210,65217,65224,65231,65237,65244,65251,65257,65264,65270,65277,65283,65289,65295,65301,65307,65313,65319,65325,65330,65336,65341,65347,65352,65357,65363,65368,65373,65378,65383,65387,65392,65397,65401,65406,65410,65415,65419,65423,65427,65431,65435,65439,65443,65447,65450,65454,65457,65461,65464,65468,65471,65474,65477,65480,65483,65486,65488,65491,65494,65496,65498,65501,65503,65505,65507,65509,65511,65513,65515,65517,65518,65520,65522,65523,65524,65526,65527,65528,65529,65530,65531,65532,65532,65533,65534,65534,65535,65535,65535,65535,65535,65535,65535,65535,65535,65535,65535,65534,65534,65533,65532,65532,65531,65530,65529,65528,65527,65526,65524,65523,65522,65520,65518,65517,65515,65513,65511,65509,65507,65505,65503,65501,65498,65496,65494,65491,65488,65486,65483,65480,65477,65474,65471,65468,65464,65461,65457,65454,65450,65447,65443,65439,65435,65431,65427,65423,65419,65415,65410,65406,65401,65397,65392,65387,65383,65378,65373,65368,65363,65357,65352,65347,65341,65336,65330,65325,65319,65313,65307,65301,65295,65289,65283,65277,65270,65264,65257,65251,65244,65237,65231,65224,65217,65210,65203,65195,65188,65181,65173,65166,65158,65151,65143,65135,65127,65119,65111,65103,65095,65087,65079,65070,65062,65053,65044,65036,65027,65018,65009,65000,64991,64982,64973,64963,64954,64944,64935,64925,64916,64906,64896,64886,64876,64866,64856,64846,64835,64825,64815,64804,64793,64783,64772,64761,64750,64739,64728,64717,64706,64695,64683,64672,64660,64649,64637,64625,64614,64602,64590,64578,64566,64553,64541,64529,64517,64504,64491,64479,64466,64453,64441,64428,64415,64402,64388,64375,64362,64349,64335,64322,64308,64294,64281,64267,64253,64239,64225,64211,64197,64182,64168,64154,64139,64125,64110,64095,64080,64066,64051,64036,64021,64005,63990,63975,63960,63944,63929,63913,63897,63882,63866,63850,63834,63818,63802,63786,63769,63753,63737,63720,63704,63687,63670,63654,63637,63620,63603,63586,63569,63552,63534,63517,63500,63482,63465,63447,63429,63412,63394,63376,63358,63340,63322,63303,63285,63267,63248,63230,63211,63193,63174,63155,63136,63118,63099,63080,63060,63041,63022,63003,62983,62964,62944,62924,62905,62885,62865,62845,62825,62805,62785,62765,62745,62724,62704,62683,62663,62642,62622,62601,62580,62559,62538,62517,62496,62475,62454,62432,62411,62389,62368,62346,62325,62303,62281,62259,62237,62215,62193,62171,62149,62127,62104,62082,62059,62037,62014,61991,61969,61946,61923,61900,61877,61854,61830,61807,61784,61761,61737,61714,61690,61666,61643,61619,61595,61571,61547,61523,61499,61475,61450,61426,61402,61377,61353,61328,61303,61279,61254,61229,61204,61179,61154,61129,61103,61078,61053,61027,61002,60976,60951,60925,60899,60874,60848,60822,60796,60770,60744,60717,60691,60665,60638,60612,60585,60559,60532,60505,60479,60452,60425,60398,60371,60344,60316,60289,60262,60234,60207,60179,60152,60124,60097,60069,60041,60013,59985,59957,59929,59901,59873,59844,59816,59788,59759,59731,59702,59673,59645,59616,59587,59558,59529,59500,59471,59442,59413,59383,59354,59325,59295,59266,59236,59206,59177,59147,59117,59087,59057,59027,58997,58967,58937,58906,58876,58845,58815,58784,58754,58723,58693,58662,58631,58600,58569,58538,58507,58476,58445,58413,58382,58351,58319,58288,58256,58225,58193,58161,58129,58098,58066,58034,58002,57969,57937,57905,57873,57841,57808,57776,57743,57711,57678,57645,57613,57580,57547,57514,57481,57448,57415,57382,57348,57315,57282,57248,57215,57182,57148,57114,57081,57047,57013,56979,56945,56912,56877,56843,56809,56775,56741,56707,56672,56638,56603,56569,56534,56500,56465,56430,56395,56361,56326,56291,56256,56221,56185,56150,56115,56080,56044,56009,55973,55938,55902,55867,55831,55795,55760,55724,55688,55652,55616,55580,55544,55508,55471,55435,55399,55362,55326,55289,55253,55216,55180,55143,55106,55069,55033,54996,54959,54922,54885,54848,54810,54773,54736,54699,54661,54624,54586,54549,54511,54474,54436,54398,54360,54323,54285,54247,54209,54171,54133,54094,54056,54018,53980,53941,53903,53865,53826,53788,53749,53710,53672,53633,53594,53555,53516,53477,53439,53399,53360,53321,53282,53243,53204,53164,53125,53086,53046,53007,52967,52927,52888,52848,52808,52769,52729,52689,52649,52609,52569,52529,52489,52449,52408,52368,52328,52287,52247,52207,52166,52126,52085,52044,52004,51963,51922,51881,51841,51800,51759,51718,51677,51636,51594,51553,51512,51471,51430,51388,51347,51305,51264,51222,51181,51139,51098,51056,51014,50972,50931,50889,50847,50805,50763,50721,50679,50637,50595,50552,50510,50468,50426,50383,50341,50298,50256,50213,50171,50128,50085,50043,50000,49957,49914,49872,49829,49786,49743,49700,49657,49614,49570,49527,49484,49441,49398,49354,49311,49267,49224,49181,49137,49093,49050,49006,48963,48919,48875,48831,48787,48744,48700,48656,48612,48568,48524,48480,48435,48391,48347,48303,48259,48214,48170,48125,48081,48037,47992,47948,47903,47858,47814,47769,47724,47680,47635,47590,47545,47500,47455,47410,47366,47320,47275,47230,47185,47140,47095,47050,47004,46959,46914,46868,46823,46778,46732,46687,46641,46596,46550,46504,46459,46413,46367,46322,46276,46230,46184,46138,46092,46046,46000,45954,45908,45862,45816,45770,45724,45678,45632,45585,45539,45493,45446,45400,45354,45307,45261,45214,45168,45121,45075,45028,44981,44935,44888,44841,44795,44748,44701,44654,44607,44561,44514,44467,44420,44373,44326,44279,44232,44184,44137,44090,44043,43996,43949,43901,43854,43807,43759,43712,43665,43617,43570,43522,43475,43427,43380,43332,43285,43237,43189,43142,43094,43046,42998,42951,42903,42855,42807,42759,42712,42664,42616,42568,42520,42472,42424,42376,42328,42280,42231,42183,42135,42087,42039,41991,41942,41894,41846,41797,41749,41701,41652,41604,41556,41507,41459,41410,41362,41313,41265,41216,41168,41119,41070,41022,40973,40924,40876,40827,40778,40729,40681,40632,40583,40534,40485,40437,40388,40339,40290,40241,40192,40143,40094,40045,39996,39947,39898,39849,39800,39751,39702,39652,39603,39554,39505,39456,39407,39357,39308,39259,39210,39160,39111,39062,39012,38963,38914,38864,38815,38765,38716,38666,38617,38568,38518,38469,38419,38370,38320,38271,38221,38171,38122,38072,38023,37973,37923,37874,37824,37774,37725,37675,37625,37576,37526,37476,37426,37377,37327,37277,37227,37177,37128,37078,37028,36978,36928,36878,36829,36779,36729,36679,36629,36579,36529,36479,36429,36379,36329,36279,36229,36179,36129,36079,36029,35979,35929,35879,35829,35779,35729,35679,35629,35579,35529,35479,35429,35379,35328,35278,35228,35178,35128,35078,35028,34978,34927,34877,34827,34777,34727,34677,34626,34576,34526,34476,34426,34375,34325,34275,34225,34175,34124,34074,34024,33974,33923,33873,33823,33773,33722,33672,33622,33572,33521,33471,33421,33371,33320,33270,33220,33170,33119,33069,33019,32969,32918,32868,32818,32768,32717,32667,32617,32566,32516,32466,32416,32365,32315,32265,32215,32164,32114,32064,32014,31963,31913,31863,31813,31762,31712,31662,31612,31561,31511,31461,31411,31360,31310,31260,31210,31160,31109,31059,31009,30959,30909,30858,30808,30758,30708,30658,30608,30557,30507,30457,30407,30357,30307,30257,30207,30156,30106,30056,30006,29956,29906,29856,29806,29756,29706,29656,29606,29556,29506,29456,29406,29356,29306,29256,29206,29156,29106,29056,29006,28956,28906,28856,28806,28756,28706,28657,28607,28557,28507,28457,28407,28358,28308,28258,28208,28158,28109,28059,28009,27959,27910,27860,27810,27761,27711,27661,27612,27562,27512,27463,27413,27364,27314,27264,27215,27165,27116,27066,27017,26967,26918,26869,26819,26770,26720,26671,26621,26572,26523,26473,26424,26375,26325,26276,26227,26178,26128,26079,26030,25981,25932,25883,25833,25784,25735,25686,25637,25588,25539,25490,25441,25392,25343,25294,25245,25196,25147,25098,25050,25001,24952,24903,24854,24806,24757,24708,24659,24611,24562,24513,24465,24416,24367,24319,24270,24222,24173,24125,24076,24028,23979,23931,23883,23834,23786,23738,23689,23641,23593,23544,23496,23448,23400,23352,23304,23255,23207,23159,23111,23063,23015,22967,22919,22871,22823,22776,22728,22680,22632,22584,22537,22489,22441,22393,22346,22298,22250,22203,22155,22108,22060,22013,21965,21918,21870,21823,21776,21728,21681,21634,21586,21539,21492,21445,21398,21351,21303,21256,21209,21162,21115,21068,21021,20974,20928,20881,20834,20787,20740,20694,20647,20600,20554,20507,20460,20414,20367,20321,20274,20228,20181,20135,20089,20042,19996,19950,19903,19857,19811,19765,19719,19673,19627,19581,19535,19489,19443,19397,19351,19305,19259,19213,19168,19122,19076,19031,18985,18939,18894,18848,18803,18757,18712,18667,18621,18576,18531,18485,18440,18395,18350,18305,18260,18215,18169,18125,18080,18035,17990,17945,17900,17855,17811,17766,17721,17677,17632,17587,17543,17498,17454,17410,17365,17321,17276,17232,17188,17144,17100,17055,17011,16967,16923,16879,16835,16791,16748,16704,16660,16616,16572,16529,16485,16442,16398,16354,16311,16268,16224,16181,16137,16094,16051,16008,15965,15921,15878,15835,15792,15749,15706,15663,15621,15578,15535,15492,15450,15407,15364,15322,15279,15237,15194,15152,15109,15067,15025,14983,14940,14898,14856,14814,14772,14730,14688,14646,14604,14563,14521,14479,14437,14396,14354,14313,14271,14230,14188,14147,14105,14064,14023,13982,13941,13899,13858,13817,13776,13735,13694,13654,13613,13572,13531,13491,13450,13409,13369,13328,13288,13248,13207,13167,13127,13086,13046,13006,12966,12926,12886,12846,12806,12766,12727,12687,12647,12608,12568,12528,12489,12449,12410,12371,12331,12292,12253,12214,12175,12136,12096,12058,12019,11980,11941,11902,11863,11825,11786,11747,11709,11670,11632,11594,11555,11517,11479,11441,11402,11364,11326,11288,11250,11212,11175,11137,11099,11061,11024,10986,10949,10911,10874,10836,10799,10762,10725,10687,10650,10613,10576,10539,10502,10466,10429,10392,10355,10319,10282,10246,10209,10173,10136,10100,10064,10027,9991,9955,9919,9883,9847,9811,9775,9740,9704,9668,9633,9597,9562,9526,9491,9455,9420,9385,9350,9314,9279,9244,9209,9174,9140,9105,9070,9035,9001,8966,8932,8897,8863,8828,8794,8760,8726,8692,8658,8623,8590,8556,8522,8488,8454,8421,8387,8353,8320,8287,8253,8220,8187,8153,8120,8087,8054,8021,7988,7955,7922,7890,7857,7824,7792,7759,7727,7694,7662,7630,7598,7566,7533,7501,7469,7437,7406,7374,7342,7310,7279,7247,7216,7184,7153,7122,7090,7059,7028,6997,6966,6935,6904,6873,6842,6812,6781,6751,6720,6690,6659,6629,6598,6568,6538,6508,6478,6448,6418,6388,6358,6329,6299,6269,6240,6210,6181,6152,6122,6093,6064,6035,6006,5977,5948,5919,5890,5862,5833,5804,5776,5747,5719,5691,5662,5634,5606,5578,5550,5522,5494,5466,5438,5411,5383,5356,5328,5301,5273,5246,5219,5191,5164,5137,5110,5083,5056,5030,5003,4976,4950,4923,4897,4870,4844,4818,4791,4765,4739,4713,4687,4661,4636,4610,4584,4559,4533,4508,4482,4457,4432,4406,4381,4356,4331,4306,4281,4256,4232,4207,4182,4158,4133,4109,4085,4060,4036,4012,3988,3964,3940,3916,3892,3869,3845,3821,3798,3774,3751,3728,3705,3681,3658,3635,3612,3589,3566,3544,3521,3498,3476,3453,3431,3408,3386,3364,3342,3320,3298,3276,3254,3232,3210,3189,3167,3146,3124,3103,3081,3060,3039,3018,2997,2976,2955,2934,2913,2893,2872,2852,2831,2811,2790,2770,2750,2730,2710,2690,2670,2650,2630,2611,2591,2571,2552,2532,2513,2494,2475,2455,2436,2417,2399,2380,2361,2342,2324,2305,2287,2268,2250,2232,2213,2195,2177,2159,2141,2123,2106,2088,2070,2053,2035,2018,2001,1983,1966,1949,1932,1915,1898,1881,1865,1848,1831,1815,1798,1782,1766,1749,1733,1717,1701,1685,1669,1653,1638,1622,1606,1591,1575,1560,1545,1530,1514,1499,1484,1469,1455,1440,1425,1410,1396,1381,1367,1353,1338,1324,1310,1296,1282,1268,1254,1241,1227,1213,1200,1186,1173,1160,1147,1133,1120,1107,1094,1082,1069,1056,1044,1031,1018,1006,994,982,969,957,945,933,921,910,898,886,875,863,852,840,829,818,807,796,785,774,763,752,742,731,720,710,700,689,679,669,659,649,639,629,619,610,600,591,581,572,562,553,544,535,526,517,508,499,491,482,473,465,456,448,440,432,424,416,408,400,392,384,377,369,362,354,347,340,332,325,318,311,304,298,291,284,278,271,265,258,252,246,240,234,228,222,216,210,205,199,194,188,183,178,172,167,162,157,152,148,143,138,134,129,125,120,116,112,108,104,100,96,92,88,85,81,78,74,71,67,64,61,58,55,52,49,47,44,41,39,37,34,32,30,28,26,24,22,20,18,17,15,13,12,11,9,8,7,6,5,4,3,3,2,1,1,0,0,0,0,0,0,0,0,0,0,0,1,1,2,3,3,4,5,6,7,8,9,11,12,13,15,17,18,20,22,24,26,28,30,32,34,37,39,41,44,47,49,52,55,58,61,64,67,71,74,78,81,85,88,92,96,100,104,108,112,116,120,125,129,134,138,143,148,152,157,162,167,172,178,183,188,194,199,205,210,216,222,228,234,240,246,252,258,265,271,278,284,291,298,304,311,318,325,332,340,347,354,362,369,377,384,392,400,408,416,424,432,440,448,456,465,473,482,491,499,508,517,526,535,544,553,562,572,581,591,600,610,619,629,639,649,659,669,679,689,700,710,720,731,742,752,763,774,785,796,807,818,829,840,852,863,875,886,898,910,921,933,945,957,969,982,994,1006,1018,1031,1044,1056,1069,1082,1094,1107,1120,1133,1147,1160,1173,1186,1200,1213,1227,1241,1254,1268,1282,1296,1310,1324,1338,1353,1367,1381,1396,1410,1425,1440,1455,1469,1484,1499,1514,1530,1545,1560,1575,1591,1606,1622,1638,1653,1669,1685,1701,1717,1733,1749,1766,1782,1798,1815,1831,1848,1865,1881,1898,1915,1932,1949,1966,1983,2001,2018,2035,2053,2070,2088,2106,2123,2141,2159,2177,2195,2213,2232,2250,2268,2287,2305,2324,2342,2361,2380,2399,2417,2436,2455,2475,2494,2513,2532,2552,2571,2591,2611,2630,2650,2670,2690,2710,2730,2750,2770,2790,2811,2831,2852,2872,2893,2913,2934,2955,2976,2997,3018,3039,3060,3081,3103,3124,3146,3167,3189,3210,3232,3254,3276,3298,3320,3342,3364,3386,3408,3431,3453,3476,3498,3521,3544,3566,3589,3612,3635,3658,3681,3705,3728,3751,3774,3798,3821,3845,3869,3892,3916,3940,3964,3988,4012,4036,4060,4085,4109,4133,4158,4182,4207,4232,4256,4281,4306,4331,4356,4381,4406,4432,4457,4482,4508,4533,4559,4584,4610,4636,4661,4687,4713,4739,4765,4791,4818,4844,4870,4897,4923,4950,4976,5003,5030,5056,5083,5110,5137,5164,5191,5219,5246,5273,5301,5328,5356,5383,5411,5438,5466,5494,5522,5550,5578,5606,5634,5662,5691,5719,5747,5776,5804,5833,5862,5890,5919,5948,5977,6006,6035,6064,6093,6122,6152,6181,6210,6240,6269,6299,6329,6358,6388,6418,6448,6478,6508,6538,6568,6598,6629,6659,6690,6720,6751,6781,6812,6842,6873,6904,6935,6966,6997,7028,7059,7090,7122,7153,7184,7216,7247,7279,7310,7342,7374,7406,7437,7469,7501,7533,7566,7598,7630,7662,7694,7727,7759,7792,7824,7857,7890,7922,7955,7988,8021,8054,8087,8120,8153,8187,8220,8253,8287,8320,8353,8387,8421,8454,8488,8522,8556,8590,8623,8658,8692,8726,8760,8794,8828,8863,8897,8932,8966,9001,9035,9070,9105,9140,9174,9209,9244,9279,9314,9350,9385,9420,9455,9491,9526,9562,9597,9633,9668,9704,9740,9775,9811,9847,9883,9919,9955,9991,10027,10064,10100,10136,10173,10209,10246,10282,10319,10355,10392,10429,10466,10502,10539,10576,10613,10650,10687,10725,10762,10799,10836,10874,10911,10949,10986,11024,11061,11099,11137,11175,11212,11250,11288,11326,11364,11402,11441,11479,11517,11555,11594,11632,11670,11709,11747,11786,11825,11863,11902,11941,11980,12019,12058,12096,12136,12175,12214,12253,12292,12331,12371,12410,12449,12489,12528,12568,12608,12647,12687,12727,12766,12806,12846,12886,12926,12966,13006,13046,13086,13127,13167,13207,13248,13288,13328,13369,13409,13450,13491,13531,13572,13613,13654,13694,13735,13776,13817,13858,13899,13941,13982,14023,14064,14105,14147,14188,14230,14271,14313,14354,14396,14437,14479,14521,14563,14604,14646,14688,14730,14772,14814,14856,14898,14940,14983,15025,15067,15109,15152,15194,15237,15279,15322,15364,15407,15450,15492,15535,15578,15621,15663,15706,15749,15792,15835,15878,15921,15965,16008,16051,16094,16137,16181,16224,16268,16311,16354,16398,16442,16485,16529,16572,16616,16660,16704,16748,16791,16835,16879,16923,16967,17011,17055,17100,17144,17188,17232,17276,17321,17365,17410,17454,17498,17543,17587,17632,17677,17721,17766,17811,17855,17900,17945,17990,18035,18080,18125,18169,18215,18260,18305,18350,18395,18440,18485,18531,18576,18621,18667,18712,18757,18803,18848,18894,18939,18985,19031,19076,19122,19168,19213,19259,19305,19351,19397,19443,19489,19535,19581,19627,19673,19719,19765,19811,19857,19903,19950,19996,20042,20089,20135,20181,20228,20274,20321,20367,20414,20460,20507,20554,20600,20647,20694,20740,20787,20834,20881,20928,20974,21021,21068,21115,21162,21209,21256,21303,21351,21398,21445,21492,21539,21586,21634,21681,21728,21776,21823,21870,21918,21965,22013,22060,22108,22155,22203,22250,22298,22346,22393,22441,22489,22537,22584,22632,22680,22728,22776,22823,22871,22919,22967,23015,23063,23111,23159,23207,23255,23304,23352,23400,23448,23496,23544,23593,23641,23689,23738,23786,23834,23883,23931,23979,24028,24076,24125,24173,24222,24270,24319,24367,24416,24465,24513,24562,24611,24659,24708,24757,24806,24854,24903,24952,25001,25050,25098,25147,25196,25245,25294,25343,25392,25441,25490,25539,25588,25637,25686,25735,25784,25833,25883,25932,25981,26030,26079,26128,26178,26227,26276,26325,26375,26424,26473,26523,26572,26621,26671,26720,26770,26819,26869,26918,26967,27017,27066,27116,27165,27215,27264,27314,27364,27413,27463,27512,27562,27612,27661,27711,27761,27810,27860,27910,27959,28009,28059,28109,28158,28208,28258,28308,28358,28407,28457,28507,28557,28607,28657,28706,28756,28806,28856,28906,28956,29006,29056,29106,29156,29206,29256,29306,29356,29406,29456,29506,29556,29606,29656,29706,29756,29806,29856,29906,29956,30006,30056,30106,30156,30207,30257,30307,30357,30407,30457,30507,30557,30608,30658,30708,30758,30808,30858,30909,30959,31009,31059,31109,31160,31210,31260,31310,31360,31411,31461,31511,31561,31612,31662,31712,31762,31813,31863,31913,31963,32014,32064,32114,32164,32215,32265,32315,32365,32416,32466,32516,32566,32617,32667,32717);
BEGIN
	Process(angle)
	variable angleCos :	integer; -- stores (90 degree - angle) to fetch cos value using sine table
	BEGIN	
		sinAngle<=sine(angle);
		angleCos := 1024-angle;					-- Calculate (90 - angle)
		if(angleCos < 0) then                   -- if result is negative add 360 degree to make it positive  
			angleCos := angleCos + 4096;
		end if;
		cosAngle <= sine(angleCos);
		--cosAngle <= sine(angle);
	end process;
	
end;

